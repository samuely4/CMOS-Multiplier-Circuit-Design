*** SPICE deck for cell HA{lay} from library Multp
*** Created on Tue Nov 13, 2018 23:17:05
*** Last revised on Sat Dec 01, 2018 12:30:47
*** Written on Sat Dec 01, 2018 12:31:02 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Multp__CR_HA FROM CELL CR_HA{lay}
.SUBCKT Multp__CR_HA A B cout gnd vdd
Mnmos@0 net@0 B gnd gnd NMOS L=0.7U W=3.5U AS=31.36P AD=13.781P PS=36.925U PD=15.75U
Mnmos@1 net@17 A gnd gnd NMOS L=0.7U W=3.5U AS=31.36P AD=11.699P PS=36.925U PD=15.05U
Mnmos@2 gnd net@17 cout gnd NMOS L=0.7U W=3.5U AS=17.191P AD=31.36P PS=25.433U PD=36.925U
Mnmos@3 cout net@0 gnd gnd NMOS L=0.7U W=3.5U AS=31.36P AD=17.191P PS=36.925U PD=25.433U
Mpmos@0 vdd B net@0 vdd PMOS L=0.7U W=7U AS=13.781P AD=47.367P PS=15.75U PD=50.167U
Mpmos@1 vdd A net@17 vdd PMOS L=0.7U W=7U AS=11.699P AD=47.367P PS=15.05U PD=50.167U
Mpmos@2 vdd net@17 net@65 vdd PMOS L=0.7U W=7U AS=10.658P AD=47.367P PS=21.35U PD=50.167U
Mpmos@3 net@65 net@0 cout vdd PMOS L=0.7U W=7U AS=17.191P AD=10.658P PS=25.433U PD=21.35U
.ENDS Multp__CR_HA

*** SUBCIRCUIT Multp__SM_HA FROM CELL SM_HA{lay}
.SUBCKT Multp__SM_HA A B gnd sum vdd
Mnmos@0 net@12 A gnd gnd NMOS L=0.7U W=3.5U AS=49.873P AD=14.7P PS=57.575U PD=16.1U
Mnmos@1 net@10 B gnd gnd NMOS L=0.7U W=3.5U AS=49.873P AD=13.781P PS=57.575U PD=15.75U
Mnmos@2 gnd net@10 net@107 gnd NMOS L=0.7U W=3.5U AS=7.074P AD=49.873P PS=14.525U PD=57.575U
Mnmos@3 net@107 net@12 sum gnd NMOS L=0.7U W=3.5U AS=9.616P AD=7.074P PS=18.9U PD=14.525U
Mnmos@4 sum A net@127 gnd NMOS L=0.7U W=3.5U AS=7.074P AD=9.616P PS=14.525U PD=18.9U
Mnmos@5 net@127 B gnd gnd NMOS L=0.7U W=3.5U AS=49.873P AD=7.074P PS=57.575U PD=14.525U
Mpmos@0 vdd A net@12 vdd PMOS L=0.7U W=7U AS=14.7P AD=51.863P PS=16.1U PD=57.225U
Mpmos@1 vdd B net@10 vdd PMOS L=0.7U W=7U AS=13.781P AD=51.863P PS=15.75U PD=57.225U
Mpmos@2 vdd net@10 net@48 vdd PMOS L=0.7U W=7U AS=19.768P AD=51.863P PS=34.563U PD=57.225U
Mpmos@3 net@48 net@12 vdd vdd PMOS L=0.7U W=7U AS=51.863P AD=19.768P PS=57.225U PD=34.563U
Mpmos@4 sum A net@48 vdd PMOS L=0.7U W=7U AS=19.768P AD=9.616P PS=34.563U PD=18.9U
Mpmos@5 net@48 B sum vdd PMOS L=0.7U W=7U AS=9.616P AD=19.768P PS=18.9U PD=34.563U
.ENDS Multp__SM_HA

*** TOP LEVEL CELL: HA{lay}
XCR_HA@0 A B cout gnd vdd Multp__CR_HA
XSM_HA@0 A B gnd sum vdd Multp__SM_HA

* Spice Code nodes in cell cell 'HA{lay}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
vA A 0 pulse(0 3.3 0 20n 40n 250n 500n)
VB B 0 pulse(0 3.3 0 20n 40n 300n 600n)
.TRANS 1.5u
.include C:\Electric\model.txt
.END
