*** SPICE deck for cell MUL{lay} from library Multp
*** Created on Tue Nov 13, 2018 23:17:36
*** Last revised on Sat Dec 01, 2018 11:23:06
*** Written on Sat Dec 01, 2018 11:23:34 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Multp__CR_FA FROM CELL CR_FA{lay}
.SUBCKT Multp__CR_FA A B cin gnd NCout vdd
Mnmos@0 net@58 A gnd gnd NMOS L=0.7U W=3.5U AS=77.338P AD=15.21P PS=87.733U PD=28.583U
Mnmos@1 gnd B net@58 gnd NMOS L=0.7U W=3.5U AS=15.21P AD=77.338P PS=28.583U PD=87.733U
Mnmos@2 net@25 B gnd gnd NMOS L=0.7U W=3.5U AS=77.338P AD=12.495P PS=87.733U PD=24.85U
Mnmos@3 NCout A net@25 gnd NMOS L=0.7U W=3.5U AS=12.495P AD=13.203P PS=24.85U PD=25.638U
Mnmos@4 net@58 cin NCout gnd NMOS L=0.7U W=3.5U AS=13.203P AD=15.21P PS=25.638U PD=28.583U
Mpmos@0 net@36 A vdd vdd PMOS L=0.7U W=7U AS=126.267P AD=15.067P PS=144.725U PD=29.75U
Mpmos@1 net@84 B net@36 vdd PMOS L=0.7U W=7U AS=15.067P AD=13.153P PS=29.75U PD=25.638U
Mpmos@2 NCout B net@84 vdd PMOS L=0.7U W=7U AS=13.153P AD=13.203P PS=25.638U PD=25.638U
Mpmos@3 net@84 A NCout vdd PMOS L=0.7U W=7U AS=13.203P AD=13.153P PS=25.638U PD=25.638U
Mpmos@4 vdd cin net@84 vdd PMOS L=0.7U W=7U AS=13.153P AD=126.267P PS=25.638U PD=144.725U
.ENDS Multp__CR_FA

*** SUBCIRCUIT Multp__SM_FA FROM CELL SM_FA{lay}
.SUBCKT Multp__SM_FA A B cin gnd NCout NSum vdd
Mnmos@0 net@84 cin gnd gnd NMOS L=0.7U W=3.5U AS=77.252P AD=9.754P PS=89.163U PD=19.162U
Mnmos@1 gnd B net@84 gnd NMOS L=0.7U W=3.5U AS=9.754P AD=77.252P PS=19.162U PD=89.163U
Mnmos@2 net@84 A gnd gnd NMOS L=0.7U W=3.5U AS=77.252P AD=9.754P PS=89.163U PD=19.162U
Mnmos@3 NSum NCout net@84 gnd NMOS L=0.7U W=3.5U AS=9.754P AD=16.678P PS=19.162U PD=30.59U
Mnmos@4 net@128 A NSum gnd NMOS L=0.7U W=3.5U AS=16.678P AD=10.841P PS=30.59U PD=21.7U
Mnmos@5 net@8 B net@128 gnd NMOS L=0.7U W=3.5U AS=10.841P AD=7.809P PS=21.7U PD=15.925U
Mnmos@6 gnd cin net@8 gnd NMOS L=0.7U W=3.5U AS=7.809P AD=77.252P PS=15.925U PD=89.163U
Mpmos@0 net@22 cin net@97 vdd PMOS L=0.7U W=7U AS=17.113P AD=13.375P PS=31.71U PD=25.725U
Mpmos@1 net@24 B net@22 vdd PMOS L=0.7U W=7U AS=13.375P AD=13.651P PS=25.725U PD=26.25U
Mpmos@2 vdd A net@24 vdd PMOS L=0.7U W=7U AS=13.651P AD=134.873P PS=26.25U PD=143.85U
Mpmos@3 net@97 NCout vdd vdd PMOS L=0.7U W=7U AS=134.873P AD=17.113P PS=143.85U PD=31.71U
Mpmos@4 NSum A net@97 vdd PMOS L=0.7U W=7U AS=17.113P AD=16.678P PS=31.71U PD=30.59U
Mpmos@5 net@97 B NSum vdd PMOS L=0.7U W=7U AS=16.678P AD=17.113P PS=30.59U PD=31.71U
Mpmos@6 NSum cin net@97 vdd PMOS L=0.7U W=7U AS=17.113P AD=16.678P PS=31.71U PD=30.59U
.ENDS Multp__SM_FA

*** SUBCIRCUIT Multp__inv_20_10 FROM CELL inv_20_10{lay}
.SUBCKT Multp__inv_20_10 gnd in out vdd
Mnmos@0 out in gnd gnd NMOS L=0.7U W=3.5U AS=19.6P AD=11.025P PS=28.7U PD=14.7U
Mpmos@0 vdd in out vdd PMOS L=0.7U W=7U AS=11.025P AD=26.95P PS=14.7U PD=35.7U
.ENDS Multp__inv_20_10

*** SUBCIRCUIT Multp__FA FROM CELL FA{lay}
.SUBCKT Multp__FA A B cin cout gnd sum vdd
XCR_FA@0 A B cin gnd net@9 vdd Multp__CR_FA
XSM_FA@0 A B cin gnd net@9 net@166 vdd Multp__SM_FA
Xinv_20_1@0 gnd net@9 cout vdd Multp__inv_20_10
Xinv_20_1@1 gnd net@166 sum vdd Multp__inv_20_10
.ENDS Multp__FA

*** SUBCIRCUIT Multp__CR_HA FROM CELL CR_HA{lay}
.SUBCKT Multp__CR_HA A B cout gnd vdd
Mnmos@0 net@0 B gnd gnd NMOS L=0.7U W=3.5U AS=31.36P AD=13.781P PS=36.925U PD=15.75U
Mnmos@1 net@17 A gnd gnd NMOS L=0.7U W=3.5U AS=31.36P AD=11.699P PS=36.925U PD=15.05U
Mnmos@2 gnd net@17 cout gnd NMOS L=0.7U W=3.5U AS=17.191P AD=31.36P PS=25.433U PD=36.925U
Mnmos@3 cout net@0 gnd gnd NMOS L=0.7U W=3.5U AS=31.36P AD=17.191P PS=36.925U PD=25.433U
Mpmos@0 vdd B net@0 vdd PMOS L=0.7U W=7U AS=13.781P AD=47.367P PS=15.75U PD=50.167U
Mpmos@1 vdd A net@17 vdd PMOS L=0.7U W=7U AS=11.699P AD=47.367P PS=15.05U PD=50.167U
Mpmos@2 vdd net@17 net@65 vdd PMOS L=0.7U W=7U AS=10.658P AD=47.367P PS=21.35U PD=50.167U
Mpmos@3 net@65 net@0 cout vdd PMOS L=0.7U W=7U AS=17.191P AD=10.658P PS=25.433U PD=21.35U
.ENDS Multp__CR_HA

*** SUBCIRCUIT Multp__SM_HA FROM CELL SM_HA{lay}
.SUBCKT Multp__SM_HA A B gnd sum vdd
Mnmos@0 net@12 A gnd gnd NMOS L=0.7U W=3.5U AS=49.873P AD=14.7P PS=57.575U PD=16.1U
Mnmos@1 net@10 B gnd gnd NMOS L=0.7U W=3.5U AS=49.873P AD=13.781P PS=57.575U PD=15.75U
Mnmos@2 gnd net@10 net@107 gnd NMOS L=0.7U W=3.5U AS=7.074P AD=49.873P PS=14.525U PD=57.575U
Mnmos@3 net@107 net@12 sum gnd NMOS L=0.7U W=3.5U AS=9.616P AD=7.074P PS=18.9U PD=14.525U
Mnmos@4 sum A net@127 gnd NMOS L=0.7U W=3.5U AS=7.074P AD=9.616P PS=14.525U PD=18.9U
Mnmos@5 net@127 B gnd gnd NMOS L=0.7U W=3.5U AS=49.873P AD=7.074P PS=57.575U PD=14.525U
Mpmos@0 vdd A net@12 vdd PMOS L=0.7U W=7U AS=14.7P AD=51.863P PS=16.1U PD=57.225U
Mpmos@1 vdd B net@10 vdd PMOS L=0.7U W=7U AS=13.781P AD=51.863P PS=15.75U PD=57.225U
Mpmos@2 vdd net@10 net@48 vdd PMOS L=0.7U W=7U AS=19.768P AD=51.863P PS=34.563U PD=57.225U
Mpmos@3 net@48 net@12 vdd vdd PMOS L=0.7U W=7U AS=51.863P AD=19.768P PS=57.225U PD=34.563U
Mpmos@4 sum A net@48 vdd PMOS L=0.7U W=7U AS=19.768P AD=9.616P PS=34.563U PD=18.9U
Mpmos@5 net@48 B sum vdd PMOS L=0.7U W=7U AS=9.616P AD=19.768P PS=18.9U PD=34.563U
.ENDS Multp__SM_HA

*** SUBCIRCUIT Multp__HA FROM CELL HA{lay}
.SUBCKT Multp__HA A B cout gnd sum vdd
XCR_HA@0 A B cout gnd vdd Multp__CR_HA
XSM_HA@0 A B gnd sum vdd Multp__SM_HA
.ENDS Multp__HA

*** SUBCIRCUIT Multp__and FROM CELL and{lay}
.SUBCKT Multp__and A AB B gnd vdd
Mnmos@0 net@7 B gnd gnd NMOS L=0.7U W=3.5U AS=27.563P AD=2.297P PS=35.175U PD=5.425U
Mnmos@1 net@1 A net@7 gnd NMOS L=0.7U W=3.5U AS=2.297P AD=9.392P PS=5.425U PD=10.5U
Mnmos@2 AB net@1 gnd gnd NMOS L=0.7U W=3.5U AS=27.563P AD=14.7P PS=35.175U PD=16.1U
Mpmos@0 net@1 B vdd vdd PMOS L=0.7U W=7U AS=30.094P AD=9.392P PS=34.44U PD=10.5U
Mpmos@1 vdd A net@1 vdd PMOS L=0.7U W=7U AS=9.392P AD=30.094P PS=10.5U PD=34.44U
Mpmos@2 AB net@1 vdd vdd PMOS L=0.7U W=7U AS=30.094P AD=14.7P PS=34.44U PD=16.1U
.ENDS Multp__and

*** TOP LEVEL CELL: MUL{lay}
XFA@1 net@515 net@518 net@505 net@529 gnd net@553 vdd Multp__FA
XFA@2 net@479 net@484 net@477 net@505 gnd net@549 vdd Multp__FA
XFA@3 net@630 net@641 net@592 net@625 gnd net@731 vdd Multp__FA
XFA@4 net@598 net@553 net@586 net@592 gnd net@588 vdd Multp__FA
XFA@5 net@657 net@556 net@625 net@684 gnd net@754 vdd Multp__FA
XFA@6 net@745 net@754 net@739 net@767 gnd out5 vdd Multp__FA
XFA@7 net@723 net@731 net@700 net@739 gnd out4 vdd Multp__FA
XFA@8 net@779 net@684 net@767 out7 gnd out6 vdd Multp__FA
XHA@3 net@465 net@461 net@477 gnd out1 vdd Multp__HA
XHA@4 net@541 net@529 net@556 gnd net@641 vdd Multp__HA
XHA@6 net@569 net@549 net@586 gnd out2 vdd Multp__HA
XHA@8 net@691 net@588 net@700 gnd out3 vdd Multp__HA
Xand@6 B1 net@541 A3 gnd vdd Multp__and
Xand@7 B1 net@515 A2 gnd vdd Multp__and
Xand@8 B1 net@479 A1 gnd vdd Multp__and
Xand@9 B1 net@465 A0 gnd vdd Multp__and
Xand@18 B0 net@518 A3 gnd vdd Multp__and
Xand@19 B0 net@484 A2 gnd vdd Multp__and
Xand@20 B0 net@461 A1 gnd vdd Multp__and
Xand@21 B0 out0 A0 gnd vdd Multp__and
Xand@22 B2 net@657 A3 gnd vdd Multp__and
Xand@23 B2 net@630 A2 gnd vdd Multp__and
Xand@24 B2 net@598 A1 gnd vdd Multp__and
Xand@25 B2 net@569 A0 gnd vdd Multp__and
Xand@26 B3 net@779 A3 gnd vdd Multp__and
Xand@27 B3 net@745 A2 gnd vdd Multp__and
Xand@28 B3 net@723 A1 gnd vdd Multp__and
Xand@29 B3 net@691 A0 gnd vdd Multp__and

* Spice Code nodes in cell cell 'MUL{lay}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
vA0 A0 0 DC 3.3
vA1 A1 0 DC 3.3
vA2 A2 0 DC 0
vA3 A3 0 DC 3.3
vB0 B0 0 DC 0
vB1 B1 0 DC 3.3
vB2 B2 0 DC 3.3
vB3 B3 0 DC 3.3
.TRANS 4u
.include C:\Electric\model.txt
.END
